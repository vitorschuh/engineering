CIRCUIT C:\Users\schuh\Desktop\f1.MSK
*
* IC Technology: K-CMOS Free-PDK-Based 45nm - 6 Metal
*
VDD 1 0 DC 1.00
V2_vdd 2 0 DC 0.20V
Vd 9 0 DC 0 PULSE(0.00 1.00 7.90N 0.10N 0.10N 7.90N 16.00N)
Vc 10 0 DC 0 PULSE(0.00 1.00 3.90N 0.10N 0.10N 3.90N 8.00N)
Vb 11 0 DC 0 PULSE(0.00 1.00 1.90N 0.10N 0.10N 1.90N 4.00N)
Va 12 0 DC 0 PULSE(0.00 1.00 0.90N 0.10N 0.10N 0.90N 2.00N)
*
* List of nodes
* "out f1" corresponds to n�3
* "N4" corresponds to n�4
* "gnd" corresponds to n�5
* "N6" corresponds to n�6
* "N7" corresponds to n�7
* "N8" corresponds to n�8
* "d" corresponds to n�9
* "c" corresponds to n�10
* "b" corresponds to n�11
* "a" corresponds to n�12
*
* MOS devices
MN1 0 4 3 0 N1  W= 0.10U L= 0.05U
MN2 6 9 4 0 N1  W= 0.40U L= 0.05U
MN3 7 10 6 0 N1  W= 0.40U L= 0.05U
MN4 8 11 7 0 N1  W= 0.40U L= 0.05U
MN5 0 12 8 0 N1  W= 0.40U L= 0.05U
MP1 2 4 3 2 P1  W= 0.10U L= 0.05U
MP2 2 9 4 2 P1  W= 0.10U L= 0.05U
MP3 4 10 2 2 P1  W= 0.10U L= 0.05U
MP4 2 11 4 2 P1  W= 0.10U L= 0.05U
MP5 4 12 2 2 P1  W= 0.10U L= 0.05U
*
C2 2 0  0.286fF
C3 3 0  0.075fF
C4 4 0  0.231fF
C6 6 0  0.082fF
C7 7 0  0.082fF
C8 8 0  0.082fF
C9 9 0  0.043fF
C10 10 0  0.040fF
C11 11 0  0.036fF
C12 12 0  0.033fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 UO=600.000 TOX= 2.0E-9
+LD =0.000U THETA=0.500 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
* (Winspice)
.options temp=27.0
.control
tran 0.1N 5.00N
print  V(11) V(10) V(9) V(2) V(5) > out.txt
plot  V(11) V(10) V(9) V(2) V(5)
.endc
.END
